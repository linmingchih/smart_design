.model Inner1_GND1_ W MODELTYPE=table N=6 RMODEL=r_Inner1_GND1_
+ LMODEL=l_Inner1_GND1_ GMODEL=g_Inner1_GND1_ CMODEL=c_Inner1_GND1_


.model r_Inner1_GND1_ sp N=6 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 15
+ 0           
+        12.11004241652989
+       0.1289579856675189
+         12.1100425893771
+       0.1289571062744238
+       0.1289578663014823
+        12.11004240637347
+       0.1289559325810503
+       0.1289568598656531
+       0.1289577288146031
+        12.11004240637348
+       0.1289548915031803
+       0.1289557342345537
+        0.128956859865662
+       0.1289578663015241
+         12.1100425893772
+       0.1289543174577367
+       0.1289548915031509
+       0.1289559325810736
+       0.1289571062745346
+       0.1289579856677385
+        12.11004241653024
+ 3162.3      
+        12.11006259958869
+       0.1289766685666422
+        12.11006432785061
+       0.1289678756376055
+       0.1289754751061833
+        12.11006249813578
+       0.1289561401900705
+       0.1289654119586986
+       0.1289741004843816
+        12.11006249813587
+       0.1289457308047765
+       0.1289541570607518
+       0.1289654119587747
+       0.1289754751065857
+        12.11006432785165
+       0.1289399911062613
+       0.1289457308045197
+       0.1289561401902772
+       0.1289678756386971
+       0.1289766685688294
+        12.11006259959215
+ 10000       
+        12.11026416903152
+       0.1291632490553851
+        12.11028143066553
+       0.1290754197220892
+       0.1291513343765502
+        12.11026316557112
+       0.1289582135239712
+       0.1290508237042634
+       0.1291376127939428
+        12.11026316557208
+       0.1288542587018263
+       0.1289384157143192
+         0.12905082370499
+        0.129151334380547
+        12.11028143067597
+        0.128796937133576
+       0.1288542586992809
+       0.1289582135260303
+       0.1290754197329469
+        0.129163249077231
+        12.11026416906615
+ 31623       
+        12.11225433419901
+        0.131004755192192
+        12.11242488264432
+       0.1301362314672417
+       0.1308875391490081
+        12.11224535016567
+       0.1289786661323886
+       0.1298942433852563
+        0.130752723160962
+        12.11224535017415
+       0.1279527127199476
+       0.1287839540325366
+       0.1298942433915033
+       0.1308875391864683
+        12.11242488274454
+       0.1273868739555328
+       0.1279527126941703
+       0.1289786661511738
+       0.1301362315720629
+       0.1310047554049381
+        12.11225433453825
+ 1e+05       
+        12.13006291383816
+       0.1474241291136387
+        12.13158820374464
+       0.1395388707335174
+       0.1463992954879521
+        12.13003896452714
+       0.1291529794882778
+        0.137436002596107
+       0.1452425100050099
+        12.13003896453229
+        0.120010481908619
+       0.1274690043215117
+       0.1374360025907206
+       0.1463992956879863
+        12.13158820444212
+       0.1149597409943941
+       0.1200104816371405
+       0.1291529795558306
+       0.1395388715045734
+       0.1474241308058593
+         12.1300629166785
+ 3.1623e+05  
+        12.23284889650019
+       0.2394146662225003
+        12.24029459494409
+       0.1895424474013885
+       0.2332447262919124
+        12.23261134266066
+       0.1290193200649078
+       0.1790018784149096
+       0.2279802124463455
+        12.23261134186786
+      0.07833367930125504
+       0.1211550842433226
+       0.1790018777369947
+       0.2332447255183672
+        12.24029459539781
+      0.05011787443630089
+      0.07833367750243211
+       0.1290193191960967
+       0.1895424489320871
+       0.2394146715271681
+        12.23284890824989
+ 1e+06       
+        12.57727429988671
+       0.5049711683090314
+        12.56895538068269
+       0.2954738400158455
+       0.4743746546681005
+        12.55453934127917
+       0.1097490565862467
+       0.2780238344065964
+       0.4717732265117127
+        12.55453934094528
+     -0.01363160039899439
+       0.1054502775234953
+       0.2780238346932841
+       0.4743746517701442
+        12.56895537226993
+     -0.08723256689639669
+     -0.01363160091808885
+       0.1097490550434134
+       0.2954738356472816
+       0.5049711641778116
+        12.57727431118156
+ 3.1623e+06  
+         13.5511966473456
+        1.017858667360179
+        13.37387164879182
+       0.3401478892679241
+       0.9391990658526161
+        13.37855323321146
+       0.0265860382150529
+       0.3662555689157074
+       0.9600240680620997
+        13.37855323848139
+     -0.08279954634302608
+       0.0693161666312718
+       0.3662555737109819
+       0.9391990681054059
+         13.3738716315511
+      -0.2142850784707586
+     -0.08279953179056299
+      0.02658604185082394
+       0.3401478675054503
+         1.01785861770875
+         13.5511966015998
+ 1e+07       
+        15.90124217432306
+        1.670070080495886
+        15.38805172489732
+       0.2180541876218536
+        1.645315926137146
+        15.40945080409736
+     -0.03902986779976592
+       0.3115556385832787
+        1.653720518210904
+        15.40945080916728
+      -0.0708554933020327
+      0.02903014716078187
+       0.3115556400357659
+        1.645315932906177
+         15.3880517234307
+      -0.3226056718914282
+     -0.07085546016967831
+      -0.0390298578880435
+        0.218054150253293
+        1.670069956026387
+        15.90124192212728
+ 3.1623e+07  
+        20.72021566303287
+        2.265776659437071
+         19.9756896042818
+      0.08413258087356335
+        2.348513046573385
+        19.97614941994039
+     -0.04902179928866657
+       0.1954037034409226
+        2.348864196905738
+        19.97614942446718
+     -0.06009809353012699
+      0.03420552331236745
+       0.1954037021617917
+        2.348513050878721
+        19.97568961870832
+      -0.3922357060659361
+     -0.06009804852579564
+     -0.04902178710014551
+      0.08413253151805497
+        2.265776445406736
+        20.72021494113835
+ 1e+08       
+        29.70421440562146
+        2.889053825167269
+         28.9256522564208
+       0.0141803772584026
+        3.045623364509841
+        28.91277833134466
+     -0.05576199884456723
+        0.132335657041029
+        3.044608530803268
+        28.91277833572811
+     -0.05860457684741041
+      0.03775368440510071
+       0.1323356545136948
+        3.045623365767631
+        28.92565226980326
+      -0.4285125623105868
+     -0.05860452585468351
+     -0.05576198687657599
+      0.01418031185695476
+        2.889053486388164
+        29.70421278933444
+ 3.1623e+08  
+         45.8982001108521
+        3.769183964291517
+        45.26018174637372
+     -0.01920991034568509
+        3.987271776629538
+        45.24444917514634
+     -0.06822653867836515
+       0.1066990087557711
+        3.986021292815649
+        45.24444917918384
+     -0.06013276892024225
+      0.03128077456245279
+        0.106699005296855
+        3.987271774167604
+          45.260181741868
+      -0.4484978543256257
+     -0.06013271502107048
+      -0.0682265290569484
+     -0.01921000188267177
+        3.769183421525641
+        45.89819687325776
+ 1e+09       
+        74.81226379026292
+        5.214612801972888
+        74.52761178850108
+     -0.03309499857067655
+         5.50780401808106
+        74.51667572825093
+     -0.08944195417460632
+       0.1034075519684707
+        5.507245775821954
+        74.51667573160562
+     -0.06461718698279187
+      0.01419819620728788
+       0.1034075475001065
+        5.507804009745145
+        74.52761174416806
+      -0.4602844795022365
+     -0.06461713198289171
+     -0.08944194978743328
+     -0.03309513520640042
+        5.214611905757163
+        74.81225765287017
+ 3.1623e+09  
+        126.2939046272297
+        7.719541123416255
+        126.6936464941742
+     -0.03351156578927439
+        8.128228836694428
+        126.6962556499748
+      -0.1262599808884342
+       0.1197479159729591
+        8.129571823450837
+        126.6962556520814
+     -0.07352650021520349
+     -0.01879647657555175
+       0.1197479100655442
+        8.128228818265955
+        126.6936463747401
+      -0.4681301533766005
+     -0.07352644548660098
+      -0.1262599864024574
+     -0.03351178183508388
+        7.719539603736861
+        126.2938933239489
+ 1e+10       
+        217.8786090470826
+         12.1375460367175
+         219.526484487915
+     -0.02084893373677099
+        12.74169931090337
+        219.5558947122421
+      -0.1911471035032544
+       0.1609796188251531
+        12.74681145255998
+        219.5558947121111
+     -0.08988713509513405
+     -0.07883872861658084
+        0.160979610557834
+        12.74169927471376
+         219.526484232569
+      -0.4747512648292707
+      -0.0898870820916689
+      -0.1911471269573253
+     -0.02084929054989296
+        12.13754341116653
+          217.87858855224
* NOTE: Solution at 1000 Hz used as DC point.

.model l_Inner1_GND1_ sp N=6 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+    3.123181131524948e-07
+    3.746976879954453e-08
+    3.101690252297039e-07
+    4.702131739618475e-09
+    3.720094855967899e-08
+    3.101353549861147e-07
+    5.904108648206075e-10
+    4.668392091956162e-09
+    3.719678658242054e-08
+    3.101353549868763e-07
+    7.414557158296325e-11
+    5.862573889380998e-10
+    4.668392092709367e-09
+    3.720094856578257e-08
+    3.101690252779272e-07
+    9.307059685575315e-12
+    7.414557208365418e-11
+    5.904108688128176e-10
+    4.702131771363737e-09
+    3.746976904891249e-08
+    3.123181140646236e-07
+ DATA = 15
+ 0           
+    6.233211456163012e-07
+    2.189461850407919e-07
+    6.092226095377317e-07
+    7.366150553560128e-08
+    2.084330301411327e-07
+     6.02294714152447e-07
+   -7.995882882180321e-09
+    6.661244768113719e-08
+    2.049691167700056e-07
+     6.02294714154177e-07
+   -6.226367783559428e-08
+   -1.158095880020408e-08
+    6.661244767959277e-08
+     2.08433030141895e-07
+     6.09222609537514e-07
+   -9.993325474541349e-08
+   -6.226367783518826e-08
+   -7.995882881767553e-09
+    7.366150553641227e-08
+    2.189461850408246e-07
+    6.233211456165601e-07
+ 3162.3      
+    6.233109458732641e-07
+    2.189364538726831e-07
+     6.09211477146238e-07
+    7.365563023269422e-08
+    2.084239217680561e-07
+    6.022846652373451e-07
+   -7.996066969407457e-09
+    6.660799731361609e-08
+    2.049608589541664e-07
+    6.022846652388359e-07
+   -6.225855158214207e-08
+   -1.157995155140322e-08
+    6.660799731186198e-08
+    2.084239217682517e-07
+    6.092114771449204e-07
+    -9.99252344055086e-08
+   -6.225855158173089e-08
+   -7.996066969383725e-09
+    7.365563023249754e-08
+     2.18936453871007e-07
+     6.23310945871182e-07
+ 10000       
+    6.232091412221075e-07
+    2.188393247128918e-07
+    6.091003586046837e-07
+    7.359698600953779e-08
+    2.083330030002967e-07
+    6.021843553401913e-07
+   -7.997907706126738e-09
+    6.656357016365349e-08
+    2.048784262060991e-07
+    6.021843553393197e-07
+   -6.220739050049408e-08
+   -1.156990479065406e-08
+    6.656357015992951e-08
+    2.083330029947726e-07
+    6.091003585923937e-07
+   -9.984518717590685e-08
+   -6.220739049980748e-08
+   -7.997907709843481e-09
+    7.359698599911538e-08
+    2.188393246939683e-07
+    6.232091411967718e-07
+ 31623       
+    6.222098882542628e-07
+    2.178858309354108e-07
+    6.080092071686571e-07
+    7.302115878403902e-08
+    2.074399155853017e-07
+    6.011987566903065e-07
+   -8.016292579977491e-09
+    6.612677836742494e-08
+    2.040683000564369e-07
+     6.01198756667174e-07
+   -6.170566156190217e-08
+   -1.147192968375828e-08
+    6.612677834520393e-08
+    2.074399155252205e-07
+    6.080092070506852e-07
+   -9.905993357511927e-08
+   -6.170566155786647e-08
+   -8.016292619133774e-09
+    7.302115867497134e-08
+    2.178858307490435e-07
+    6.222098880022384e-07
+ 1e+05       
+    6.137214601028567e-07
+    2.097780314353127e-07
+    5.987090582214253e-07
+    6.811734805048378e-08
+    1.998091880036646e-07
+    5.927592695997705e-07
+   -8.192546488173405e-09
+    6.236966064315432e-08
+    1.971196999119371e-07
+    5.927592694467811e-07
+   -5.747394503828021e-08
+   -1.068192968323328e-08
+    6.236966051691569e-08
+     1.99809187584398e-07
+     5.98709057340661e-07
+   -9.242170371360317e-08
+   -5.747394496573312e-08
+   -8.192546746219771e-09
+    6.811734721898236e-08
+    2.097780299536965e-07
+    6.137214580308107e-07
+ 3.1623e+05  
+    5.767530875021992e-07
+    1.744596768418505e-07
+    5.578943707728587e-07
+    4.681470707244658e-08
+    1.661401725674966e-07
+    5.551581718684977e-07
+    -9.11768616669513e-09
+    4.551825993043168e-08
+    1.660327429167678e-07
+    5.551581718739397e-07
+   -3.963159347984779e-08
+   -7.825424733841379e-09
+    4.551825998161765e-08
+    1.661401719327388e-07
+    5.578943684921908e-07
+   -6.432033767664282e-08
+   -3.963159266301437e-08
+   -9.117686368896764e-09
+    4.681470469322903e-08
+    1.744596716994722e-07
+    5.767530793418466e-07
+ 1e+06       
+    5.177705392710746e-07
+    1.202149170854461e-07
+    4.948402955753534e-07
+    1.683610315004872e-08
+    1.150424511323277e-07
+    4.956358500587726e-07
+   -9.019221978178819e-09
+    2.049691007356099e-08
+    1.170864312541967e-07
+    4.956358505979426e-07
+   -1.491474512736322e-08
+    -4.34272358670092e-09
+    2.049691052603831e-08
+    1.150424513834913e-07
+    4.948402942429045e-07
+   -2.631159535747494e-08
+   -1.491474341983825e-08
+   -9.019221503996522e-09
+    1.683610083993244e-08
+    1.202149107395772e-07
+    5.177705268068414e-07
+ 3.1623e+06  
+    4.579267827848218e-07
+    7.566640557863115e-08
+    4.407381521790768e-07
+    2.360498931898909e-09
+    7.583192544509456e-08
+    4.417078434608743e-07
+   -3.909263502363222e-09
+    5.643811214661851e-09
+      7.6144702983869e-08
+    4.417078436127794e-07
+   -1.825400688506183e-09
+   -1.724485004636418e-09
+    5.643811235241337e-09
+    7.583192572130883e-08
+    4.407381524138287e-07
+   -7.451498592603879e-09
+   -1.825399674247334e-09
+   -3.909263167943773e-09
+    2.360497901643459e-09
+    7.566640163566612e-08
+    4.579267713087721e-07
+ 1e+07       
+    4.050934593833404e-07
+    5.093607385090749e-08
+    3.978085249908725e-07
+    2.402582464148626e-09
+     5.22460765214613e-08
+    3.977031714108724e-07
+   -1.616561452759447e-10
+    3.151936481448903e-09
+    5.207541553914121e-08
+    3.977031714097713e-07
+    1.342813295493764e-10
+    2.495363688032402e-10
+    3.151936430560214e-09
+    5.224607653658522e-08
+    3.978085252927371e-07
+   -1.879934366687063e-09
+    1.342816258321075e-10
+   -1.616560649977478e-10
+     2.40258218595661e-09
+    5.093607222549092e-08
+    4.050934514435431e-07
+ 3.1623e+07  
+    3.663958181542891e-07
+    4.196350092534995e-08
+    3.635200647882617e-07
+    4.096754690054378e-09
+    4.224546018721777e-08
+    3.634029765973108e-07
+    4.888486154136909e-10
+    4.171127131304086e-09
+    4.221721260307053e-08
+    3.634029765970913e-07
+    8.987268647014259e-11
+    5.789684912244213e-10
+    4.171127120330787e-09
+    4.224546017779388e-08
+    3.635200648613888e-07
+   -3.665695562546919e-10
+    8.987274762015872e-11
+    4.888486259923775e-10
+    4.096754611058833e-09
+    4.196350036169641e-08
+    3.663958137213126e-07
+ 1e+08       
+    3.419633816247335e-07
+    3.924664670295258e-08
+    3.399432247073794e-07
+     4.58745861225851e-09
+    3.912844087351525e-08
+    3.398956773689571e-07
+    5.619151775849235e-10
+    4.575975533536986e-09
+     3.91215841334511e-08
+    3.398956773691231e-07
+     7.34634228976146e-11
+    5.768068874645407e-10
+    4.575975531686753e-09
+     3.91284408723791e-08
+    3.399432247320445e-07
+   -6.002099682314485e-11
+     7.34634341378117e-11
+    5.619151787936595e-10
+     4.58745859371667e-09
+    3.924664656483868e-08
+    3.419633795761027e-07
+ 3.1623e+08  
+    3.276593838862505e-07
+    3.827008742999618e-08
+    3.256712989982506e-07
+    4.683332672591657e-09
+     3.80495222774292e-08
+    3.256380026805407e-07
+    5.784305775835939e-10
+    4.656466882135611e-09
+    3.804535224545795e-08
+    3.256380026809526e-07
+    7.220738602356179e-11
+    5.781545565800131e-10
+    4.656466882176373e-09
+    3.804952228027276e-08
+    3.256712990273092e-07
+    -3.41814285001914e-12
+    7.220738819635575e-11
+    5.784305790898304e-10
+    4.683332679953298e-09
+    3.827008748898731e-08
+    3.276593832611948e-07
+ 1e+09       
+    3.195104809470625e-07
+    3.782633308024827e-08
+    3.174517355451731e-07
+    4.699777858331245e-09
+    3.757535179359358e-08
+    3.174195050112641e-07
+     5.85146672231803e-10
+    4.668606972448912e-09
+    3.757138564326096e-08
+     3.17419505011854e-07
+    7.298881967671813e-11
+    5.818637190449119e-10
+    4.668606972966326e-09
+    3.757535179825573e-08
+    3.174517355832995e-07
+    6.937794924344568e-12
+    7.298882035449218e-11
+    5.851466748976192e-10
+    4.699777878894324e-09
+    3.782633324195089e-08
+    3.195104811377507e-07
+ 3.1623e+09  
+      3.1490906392387e-07
+    3.759591842012852e-08
+    3.127943561401773e-07
+    4.702084186336632e-09
+    3.733292968988733e-08
+     3.12761363333616e-07
+    5.885550385180286e-10
+    4.669191920983004e-09
+     3.73288622616824e-08
+    3.127613633343148e-07
+    7.369824074366973e-11
+    5.845979944324558e-10
+    4.669191921663338e-09
+    3.733292969548277e-08
+    3.127943561846256e-07
+    8.895904309564339e-12
+    7.369824123340069e-11
+    5.885550420126885e-10
+    4.702084214084151e-09
+    3.759591863811201e-08
+    3.149090645760153e-07
+ 1e+10       
+    3.123181131524948e-07
+    3.746976879954453e-08
+    3.101690252297039e-07
+    4.702131739618475e-09
+    3.720094855967899e-08
+    3.101353549861147e-07
+    5.904108648206075e-10
+    4.668392091956162e-09
+    3.719678658242054e-08
+    3.101353549868763e-07
+    7.414557158296325e-11
+    5.862573889380998e-10
+    4.668392092709367e-09
+    3.720094856578257e-08
+    3.101690252779272e-07
+    9.307059685575315e-12
+    7.414557208365418e-11
+    5.904108688128176e-10
+    4.702131771363737e-09
+    3.746976904891249e-08
+    3.123181140646236e-07
* NOTE: Solution at 1000 Hz used as DC point.

.model g_Inner1_GND1_ sp N=6 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ DATA = 15
+ 0           
+    8.643921080237854e-11
+   -1.055154279185852e-11
+     8.83423139947805e-11
+    -5.59777185192315e-14
+   -1.054163471118698e-11
+    8.834236569860033e-11
+     -2.6496079833565e-16
+   -5.592384668220514e-14
+    -1.05416344298984e-11
+      8.8342365698599e-11
+    1.052563486753266e-16
+   -2.768614846776194e-16
+      -5.592384676288e-14
+   -1.054163471126151e-11
+    8.834231399403092e-11
+    1.196632386913854e-16
+    1.052514172197475e-16
+   -2.649662016875797e-16
+   -5.597772459210375e-14
+   -1.055154286154011e-11
+    8.643920541299805e-11
+ 3162.3      
+    8.620002095559643e-10
+   -1.052304852817119e-10
+    8.809812973383834e-10
+   -5.581642297903733e-13
+   -1.051316822409189e-10
+    8.809818128279941e-10
+   -2.644591888259051e-15
+     -5.5762676989261e-13
+   -1.051316794350179e-10
+    8.809818128279816e-10
+    9.748846722852183e-16
+   -2.762892933974735e-15
+   -5.576267707011179e-13
+   -1.051316822416613e-10
+    8.809812973308916e-10
+    1.107889310357032e-15
+    9.748392100333562e-16
+   -2.644646030527042e-15
+   -5.581642904023953e-13
+   -1.052304859797392e-10
+    8.620001551146272e-10
+ 10000       
+    8.422708429456899e-09
+   -1.028365573643424e-09
+    8.608231252855443e-09
+   -5.452570754471623e-12
+   -1.027400231027768e-09
+      8.6082362873321e-09
+   -2.589468965372694e-14
+   -5.447313663911602e-12
+    -1.02740020359061e-09
+    8.608236287331978e-09
+    1.098031604079241e-14
+   -2.704217447208841e-14
+   -5.447313671892071e-12
+   -1.027400231034998e-09
+    8.608231252781898e-09
+    1.250903671540988e-14
+    1.097978893679245e-14
+   -2.589522388969279e-14
+   -5.452571347569524e-12
+   -1.028365580528588e-09
+    8.422707883087384e-09
+ 31623       
+    6.902389084068925e-08
+   -8.439163799693786e-09
+    7.054877876077156e-08
+   -4.457690124388893e-11
+   -8.431258844990326e-09
+    7.054881982147817e-08
+   -2.159929329297315e-13
+   -4.453344081396948e-11
+   -8.431258618858607e-09
+    7.054881982147723e-08
+    -6.48341299600174e-14
+   -2.247766242211931e-13
+   -4.453344088606158e-11
+   -8.431258845047987e-09
+    7.054877876014053e-08
+   -7.460893058747964e-14
+   -6.483064871450891e-14
+   -2.159977436188769e-13
+   -4.457690619264339e-11
+   -8.439163861359462e-09
+    6.902388520087721e-08
+ 1e+05       
+    3.212279696705432e-07
+   -3.934056777839199e-08
+    3.283500157861708e-07
+   -2.068362839516134e-10
+   -3.930381490012775e-08
+    3.283502057487498e-07
+   -1.006990266589134e-12
+   -2.066341176806703e-10
+   -3.930381385271808e-08
+    3.283502057487453e-07
+   -3.475114992955428e-13
+   -1.046462412412586e-12
+   -2.066341180612509e-10
+   -3.930381490039799e-08
+    3.283500157830436e-07
+   -4.030202170944003e-13
+   -3.474911542369463e-13
+   -1.007015551500271e-12
+   -2.068363081620656e-10
+   -3.934056809607644e-08
+    3.212279368384818e-07
+ 3.1623e+05  
+    1.233969828603122e-06
+   -1.512343942451716e-07
+    1.261371395392203e-06
+   -7.934673207870338e-10
+   -1.510932749350444e-07
+    1.261372123172083e-06
+   -3.837702947094935e-12
+   -7.926946973320117e-10
+   -1.510932709409557e-07
+    1.261372123172065e-06
+   -1.344183880993646e-12
+   -3.990535611890249e-12
+   -7.926946988829344e-10
+   -1.510932749361043e-07
+    1.261371395379814e-06
+   -1.563220880080132e-12
+    -1.34410255304996e-12
+   -3.837805761952368e-12
+    -7.93467416946586e-10
+    -1.51234395519494e-07
+    1.233969691270906e-06
+ 1e+06       
+     4.35687524624628e-06
+    -5.34164604555158e-07
+    4.453697156028241e-06
+    -2.79959961626959e-09
+   -5.336664647980309e-07
+     4.45369972218498e-06
+     -1.3377053865611e-11
+   -2.796892212652836e-09
+   -5.336664508218464e-07
+    4.453699722184915e-06
+   -4.875567606784755e-12
+   -1.393159009611742e-11
+   -2.796892218327279e-09
+   -5.336664648018775e-07
+    4.453697155983664e-06
+   -5.668797807201832e-12
+   -4.875271581734305e-12
+   -1.337742946492155e-11
+   -2.799599965373501e-09
+   -5.341646091545441e-07
+    4.356874741831533e-06
+ 3.1623e+06  
+    1.460088969932716e-05
+   -1.790413498318545e-06
+    1.492547963884455e-05
+   -9.378467766767774e-09
+   -1.788744362854512e-06
+    1.492548823241935e-05
+   -4.407693024620897e-11
+   -9.369481725685014e-09
+   -1.788744316517509e-06
+    1.492548823241913e-05
+   -1.699384821369585e-11
+   -4.600976518834406e-11
+   -9.369481745204349e-09
+   -1.788744362867834e-06
+    1.492547963869304e-05
+   -1.972316465236527e-11
+   -1.699282832273765e-11
+   -4.407822053492485e-11
+   -9.378468968582658e-09
+   -1.790413513924582e-06
+    1.460088797588319e-05
+ 1e+07       
+    4.723916640976657e-05
+   -5.793011236462051e-06
+    4.828947576952002e-05
+   -3.033623035443879e-08
+    -5.78761149288393e-06
+    4.828950356261856e-05
+   -1.396470006283993e-10
+   -3.030749577499938e-08
+   -5.787611344857379e-06
+     4.82895035626178e-05
+   -5.769916625019675e-11
+   -1.462082281139448e-10
+   -3.030749583955483e-08
+   -5.787611492928683e-06
+    4.828947576902392e-05
+   -6.678414040988533e-11
+   -5.769577428393301e-11
+   -1.396512623484495e-10
+    -3.03362343523765e-08
+   -5.793011287323391e-06
+    4.723916078652017e-05
+ 3.1623e+07  
+    0.0001491890480441925
+   -1.829526258254165e-05
+    0.0001525060847854306
+   -9.579598904729663e-08
+   -1.827821043842123e-05
+    0.0001525061725469381
+   -4.301025960284245e-10
+   -9.570648450424929e-08
+   -1.827820997778307e-05
+    0.0001525061725469356
+   -1.925097977952799e-10
+   -4.519868267634578e-10
+   -9.570648471233263e-08
+   -1.827821043856862e-05
+    0.0001525060847838462
+   -2.221005205660199e-10
+   -1.924987741544259e-10
+   -4.301163141605222e-10
+   -9.579600205134481e-08
+   -1.829526274387931e-05
+    0.0001491890302510069
+ 1e+08       
+     0.000463953958467721
+    -5.68930502913708e-05
+    0.0004742685112214681
+   -2.978930457170757e-07
+   -5.684002363254264e-05
+    0.0004742687841356843
+   -1.299229573594853e-09
+    -2.97619053698492e-07
+   -5.684002222387218e-05
+    0.0004742687841356762
+   -6.351416586944107e-10
+   -1.371404787597211e-09
+   -2.976190543588123e-07
+   -5.684002363302213e-05
+    0.0004742685112164855
+   -7.302507713973585e-10
+   -6.351063327867367e-10
+   -1.299273042678723e-09
+   -2.978930874389604e-07
+    -5.68930507945547e-05
+    0.0004639539032356717
+ 3.1623e+08  
+     0.001432507525155634
+   -0.0001756537837633322
+     0.001464351038705384
+   -9.197393165904756e-07
+    -0.000175490066343029
+     0.001464351881359356
+   -3.884353453578276e-09
+   -9.189077691784424e-07
+   -0.0001754900620725484
+     0.001464351881359329
+   -2.082435801973657e-09
+   -4.120905306725809e-09
+   -9.189077712596623e-07
+   -0.0001754900663445793
+     0.001464351038689822
+   -2.386274914513803e-09
+   -2.082323314640473e-09
+   -3.884490251716497e-09
+   -9.197394496143961e-07
+   -0.0001756537853208045
+     0.001432507355164208
+ 1e+09       
+     0.004429879781128581
+   -0.0005431680102143139
+     0.004528343453397979
+   -2.844019241581988e-06
+   -0.0005426617597621944
+     0.004528346059108659
+   -1.161929536330724e-08
+   -2.841492356744691e-06
+   -0.0005426617468006652
+     0.004528346059108573
+   -6.813322031841978e-09
+   -1.239299089586537e-08
+   -2.841492363316204e-06
+    -0.000542661759767205
+     0.004528343453349285
+   -7.784535667826472e-09
+   -6.812963525677424e-09
+   -1.161972664276271e-08
+   -2.844019666005868e-06
+   -0.0005431680150455652
+     0.004429879256456084
+ 3.1623e+09  
+      0.01385073269098723
+    -0.001698303851830762
+      0.01415859527841314
+   -8.891177094441803e-06
+    -0.001696721092736025
+      0.01415860342416793
+   -3.524327203996284e-08
+   -8.883399994008045e-06
+    -0.001696721052892572
+      0.01415860342416765
+   -2.232510744662527e-08
+   -3.777782084543129e-08
+   -8.883400014974953e-06
+    -0.001696721092752291
+      0.01415859527825914
+   -2.545113404959994e-08
+   -2.232395585341435e-08
+    -3.52446460925222e-08
+   -8.891178458633718e-06
+    -0.001698303867007978
+      0.01385073104678786
+ 1e+10       
+      0.04421072934111418
+      -0.0054212891340467
+      0.04519356292083585
+   -2.837386748809331e-05
+    -0.005416237534517599
+       0.0451935889115602
+   -1.100515342328646e-07
+   -2.834932302416158e-05
+    -0.005416237408914347
+      0.04519358891155927
+    -7.34888749899721e-08
+   -1.183937747708932e-07
+   -2.834932309230731e-05
+    -0.005416237534570883
+      0.04519356292033914
+   -8.367954744216674e-08
+   -7.348512267344379e-08
+   -1.100559948478571e-07
+   -2.837387193262945e-05
+    -0.005421289182837912
+      0.04421072404460569
* NOTE: Solution at 1000 Hz used as DC point.

.model c_Inner1_GND1_ sp N=6 SPACING=nonuniform VALTYPE=real
+ INTERPOLATION=spline
+ INFINITY =
+    1.304558178558076e-10
+   -1.573137465881948e-11
+    1.332533638392311e-10
+   -8.623305321665502e-14
+   -1.571632315426767e-11
+    1.332534451007411e-10
+   -3.292967321970928e-16
+   -8.615892329894515e-14
+   -1.571632275605218e-11
+    1.332534451007384e-10
+    2.592825155504884e-16
+    -3.58343164184975e-16
+   -8.615892331367102e-14
+   -1.571632315441083e-11
+    1.332533638385529e-10
+    2.811198840215994e-16
+    2.592770341376118e-16
+   -3.292979610091551e-16
+   -8.623306121740331e-14
+   -1.573137467820262e-11
+    1.304558288372686e-10
+ DATA = 15
+ 0           
+    1.363309704085514e-10
+   -1.645155354975559e-11
+    1.392590276808433e-10
+   -9.000841302744904e-14
+    -1.64358303546622e-11
+    1.392591124036402e-10
+    -3.46270299070088e-16
+   -8.993075290960633e-14
+   -1.643582993825657e-11
+    1.392591124036373e-10
+    2.668825515529862e-16
+   -3.761802311580891e-16
+   -8.993075293230441e-14
+   -1.643583035481113e-11
+    1.392590276801037e-10
+    2.898733686261049e-16
+    2.668766433444976e-16
+   -3.462720538047356e-16
+   -9.000842153328102e-14
+   -1.645155357534965e-11
+     1.36330980719395e-10
+ 3162.3      
+    1.363288346196866e-10
+   -1.645129381943295e-11
+    1.392568452488562e-10
+   -9.000702093763565e-14
+   -1.643557086965849e-11
+    1.392569299703589e-10
+   -3.462640572635479e-16
+   -8.992936212055543e-14
+   -1.643557045325972e-11
+     1.39256929970356e-10
+     2.66879491190681e-16
+   -3.761736447012767e-16
+   -8.992936214325192e-14
+   -1.643557086980744e-11
+    1.392568452481164e-10
+    2.898699565752445e-16
+    2.668735830929365e-16
+   -3.462658119013045e-16
+   -9.000702944332578e-14
+   -1.645129384502571e-11
+    1.363288449305658e-10
+ 10000       
+    1.363124608892484e-10
+   -1.644930426355665e-11
+    1.392401145654384e-10
+    -8.99963339136534e-14
+     -1.6433583195312e-11
+    1.392401992769933e-10
+   -3.462168103883532e-16
+   -8.991868500709062e-14
+   -1.643358277896552e-11
+    1.392401992769906e-10
+    2.668551700643134e-16
+   -3.761236607910519e-16
+   -8.991868502977716e-14
+   -1.643358319546093e-11
+    1.392401145646988e-10
+    2.898429353640074e-16
+    2.668492627958064e-16
+   -3.462185643408378e-16
+   -8.999634241826277e-14
+   -1.644930428914033e-11
+    1.363124712002403e-10
+ 31623       
+    1.361824699220171e-10
+   -1.643346281727598e-11
+    1.391072718336229e-10
+   -8.991190907766214e-14
+   -1.641775666303069e-11
+    1.391073564669771e-10
+   -3.458241236425949e-16
+   -8.983434064692415e-14
+   -1.641775624710605e-11
+    1.391073564669743e-10
+    2.666868015847573e-16
+   -3.757119747464138e-16
+   -8.983434066950564e-14
+    -1.64177566631795e-11
+    1.391072718328844e-10
+    2.896532078748652e-16
+    2.666809013521592e-16
+   -3.458258705094529e-16
+   -8.991191757343445e-14
+   -1.643346284276683e-11
+     1.36182480238488e-10
+ 1e+05       
+    1.357330194602863e-10
+   -1.637841281799062e-11
+    1.386478540828181e-10
+   -8.962252626864879e-14
+   -1.636275808813724e-11
+    1.386479384504345e-10
+   -3.443727822023273e-16
+   -8.954524550583567e-14
+   -1.636275767370409e-11
+    1.386479384504317e-10
+    2.662415557713881e-16
+   -3.742100331020097e-16
+   -8.954524552789674e-14
+    -1.63627580882857e-11
+     1.38647854082084e-10
+    2.891336103203591e-16
+     2.66235682906316e-16
+   -3.443744944403433e-16
+   -8.962253473192081e-14
+   -1.637841284303694e-11
+    1.357330298231671e-10
+ 3.1623e+05  
+    1.352445740315184e-10
+   -1.631855638507451e-11
+    1.381485649341757e-10
+   -8.930834916131442e-14
+   -1.630295752184994e-11
+    1.381486490135532e-10
+   -3.428235259210049e-16
+     -8.9231377697259e-14
+   -1.630295710901733e-11
+    1.381486490135504e-10
+    2.657366361730167e-16
+   -3.726033622284888e-16
+   -8.923137771872266e-14
+   -1.630295752199799e-11
+    1.381485649334464e-10
+    2.885446842341051e-16
+    2.657307944847984e-16
+   -3.428251985016981e-16
+   -8.930835758771285e-14
+   -1.631855640962172e-11
+    1.352445844479533e-10
+ 1e+06       
+    1.347386953095319e-10
+   -1.625654829414853e-11
+    1.376314495739613e-10
+    -8.89831363810934e-14
+   -1.624100727967144e-11
+    1.376315333551178e-10
+   -3.412523323245592e-16
+   -8.890648138551817e-14
+   -1.624100686847419e-11
+    1.376315333551149e-10
+    2.651849901685897e-16
+   -3.709694359553126e-16
+   -8.890648140633963e-14
+   -1.624100727981906e-11
+    1.376314495732371e-10
+     2.87902831315097e-16
+    2.651791820472975e-16
+   -3.412539623484576e-16
+   -8.898314476784645e-14
+   -1.625654831816944e-11
+    1.347387057830739e-10
+ 3.1623e+06  
+    1.342186478849772e-10
+   -1.619279146838298e-11
+    1.370998461752047e-10
+   -8.864896212216281e-14
+   -1.617730991280266e-11
+     1.37099929650037e-10
+   -3.396708988462278e-16
+   -8.857262855829041e-14
+   -1.617730950326428e-11
+    1.370999296500341e-10
+    2.645882247917348e-16
+   -3.693201403891701e-16
+    -8.85726285784303e-14
+   -1.617730991294981e-11
+    1.370998461744858e-10
+    2.872101952469823e-16
+    2.645824523951944e-16
+   -3.396724837773889e-16
+   -8.864897046675658e-14
+     -1.6192791491855e-11
+    1.342186584185388e-10
+ 1e+07       
+    1.336876963485044e-10
+   -1.612768883094812e-11
+    1.365570929109358e-10
+   -8.830790057869972e-14
+   -1.611226797244447e-11
+    1.365571760732196e-10
+   -3.380909229192489e-16
+   -8.823189120325289e-14
+   -1.611226756457721e-11
+    1.365571760732167e-10
+    2.639479470760795e-16
+     -3.6766736163675e-16
+    -8.82318912226773e-14
+   -1.611226797259113e-11
+    1.365570929102224e-10
+    2.864689197134088e-16
+    2.639422123298699e-16
+   -3.380924605852592e-16
+   -8.830790887887813e-14
+   -1.612768885385326e-11
+     1.33687706944358e-10
+ 3.1623e+07  
+     1.33149105290764e-10
+   -1.606164330501425e-11
+    1.360065279541842e-10
+    -8.79620259448812e-14
+   -1.604628400979777e-11
+    1.360066107995744e-10
+   -3.365241019768601e-16
+   -8.788634130808279e-14
+   -1.604628360360258e-11
+    1.360066107995716e-10
+    2.632657640552515e-16
+   -3.660229858047411e-16
+   -8.788634132676329e-14
+    -1.60462840099439e-11
+    1.360065279534765e-10
+    2.856811483980241e-16
+    2.632600686527052e-16
+   -3.365255905688355e-16
+   -8.796203419864603e-14
+    -1.60616433273391e-11
+    1.331491159505414e-10
+ 1e+08       
+    1.326061393024063e-10
+   -1.599505781375164e-11
+    1.354514894779799e-10
+   -8.761341241488436e-14
+   -1.597976057606344e-11
+    1.354515720040104e-10
+   -3.349821334522994e-16
+   -8.753805086045731e-14
+   -1.597976017152999e-11
+    1.354515720040076e-10
+    2.625432827628784e-16
+   -3.643988989998324e-16
+   -8.753805087837093e-14
+   -1.597976057620902e-11
+    1.354514894772781e-10
+    2.848490249844758e-16
+    2.625376281650811e-16
+    -3.34983571524885e-16
+   -8.761342062049524e-14
+    -1.59950578354874e-11
+    1.326061500270988e-10
+ 3.1623e+08  
+    1.320620629740815e-10
+   -1.592833528033058e-11
+    1.348953156553526e-10
+   -8.726413418288624e-14
+   -1.591310022244238e-11
+    1.348953978614362e-10
+   -3.334767147788044e-16
+   -8.718909184805362e-14
+   -1.591309981954905e-11
+    1.348953978614334e-10
+    2.617821102325879e-16
+   -3.628069873287127e-16
+   -8.718909186518287e-14
+   -1.591310022258738e-11
+    1.348953156546567e-10
+    2.839746931564116e-16
+    2.617764976683788e-16
+   -3.334781012501746e-16
+   -8.726414233886065e-14
+   -1.592833530147302e-11
+    1.320620737640403e-10
+ 1e+09       
+    1.315201408964399e-10
+   -1.586187862792134e-11
+    1.343413446593322e-10
+   -8.691626544306394e-14
+   -1.584670550013547e-11
+    1.343414265467607e-10
+   -3.320195433896131e-16
+   -8.684153625854892e-14
+   -1.584670509884937e-11
+     1.34341426546758e-10
+    2.609838534980077e-16
+   -3.612591368980706e-16
+   -8.684153627488176e-14
+   -1.584670550027988e-11
+    1.343413446586422e-10
+    2.830602965974789e-16
+    2.609782839639792e-16
+   -3.320208775414714e-16
+   -8.691627354817718e-14
+   -1.586187864847085e-11
+    1.315201517513759e-10
+ 3.1623e+09  
+    1.309836376601318e-10
+   -1.579609077969422e-11
+    1.337929146629485e-10
+    -8.65718803895945e-14
+   -1.578097896034361e-11
+    1.337929962348928e-10
+   -3.306223167179633e-16
+   -8.649745607962038e-14
+   -1.578097856062054e-11
+      1.3379299623489e-10
+    2.601501195927653e-16
+   -3.597672338145951e-16
+   -8.649745609515026e-14
+    -1.57809789604874e-11
+    1.337929146622644e-10
+    2.821079789913256e-16
+    2.601445938532632e-16
+   -3.306235981955425e-16
+   -8.657188844287977e-14
+   -1.579609079965576e-11
+    1.309836485791153e-10
+ 1e+10       
+    1.304558178558076e-10
+   -1.573137465881948e-11
+    1.332533638392311e-10
+   -8.623305321665502e-14
+   -1.571632315426767e-11
+    1.332534451007411e-10
+   -3.292967321970928e-16
+   -8.615892329894515e-14
+   -1.571632275605218e-11
+    1.332534451007384e-10
+    2.592825155504884e-16
+    -3.58343164184975e-16
+   -8.615892331367102e-14
+   -1.571632315441083e-11
+    1.332533638385529e-10
+    2.811198840215994e-16
+    2.592770341376118e-16
+   -3.292979610091551e-16
+   -8.623306121740331e-14
+   -1.573137467820262e-11
+    1.304558288372686e-10
* NOTE: Solution at 1000 Hz used as DC point.

